`timescale 1ns / 1ps

module carry_save_adder(
    input [63:0] sayi1, sayi2,
    output [63:0] toplam
    );

    wire [63:0] carry1, carry2, sum;

    full_adder fa_1_1(sayi1[0], sayi2[0], 1'b0, sum[0], carry1[0]);
    full_adder fa_1_2(sayi1[1], sayi2[1], 1'b0, sum[1], carry1[1]);
    full_adder fa_1_3(sayi1[2], sayi2[2], 1'b0, sum[2], carry1[2]);
    full_adder fa_1_4(sayi1[3], sayi2[3], 1'b0, sum[3], carry1[3]);
    full_adder fa_1_5(sayi1[4], sayi2[4], 1'b0, sum[4], carry1[4]);
    full_adder fa_1_6(sayi1[5], sayi2[5], 1'b0, sum[5], carry1[5]);
    full_adder fa_1_7(sayi1[6], sayi2[6], 1'b0, sum[6], carry1[6]);
    full_adder fa_1_8(sayi1[7], sayi2[7], 1'b0, sum[7], carry1[7]);
    full_adder fa_1_9(sayi1[8], sayi2[8], 1'b0, sum[8], carry1[8]);
    full_adder fa_1_10(sayi1[9], sayi2[9], 1'b0, sum[9], carry1[9]);
    full_adder fa_1_11(sayi1[10], sayi2[10], 1'b0, sum[10], carry1[10]);
    full_adder fa_1_12(sayi1[11], sayi2[11], 1'b0, sum[11], carry1[11]);
    full_adder fa_1_13(sayi1[12], sayi2[12], 1'b0, sum[12], carry1[12]);
    full_adder fa_1_14(sayi1[13], sayi2[13], 1'b0, sum[13], carry1[13]);
    full_adder fa_1_15(sayi1[14], sayi2[14], 1'b0, sum[14], carry1[14]);
    full_adder fa_1_16(sayi1[15], sayi2[15], 1'b0, sum[15], carry1[15]);
    full_adder fa_1_17(sayi1[16], sayi2[16], 1'b0, sum[16], carry1[16]);
    full_adder fa_1_18(sayi1[17], sayi2[17], 1'b0, sum[17], carry1[17]);
    full_adder fa_1_19(sayi1[18], sayi2[18], 1'b0, sum[18], carry1[18]);
    full_adder fa_1_20(sayi1[19], sayi2[19], 1'b0, sum[19], carry1[19]);
    full_adder fa_1_21(sayi1[20], sayi2[20], 1'b0, sum[20], carry1[20]);
    full_adder fa_1_22(sayi1[21], sayi2[21], 1'b0, sum[21], carry1[21]);
    full_adder fa_1_23(sayi1[22], sayi2[22], 1'b0, sum[22], carry1[22]);
    full_adder fa_1_24(sayi1[23], sayi2[23], 1'b0, sum[23], carry1[23]);
    full_adder fa_1_25(sayi1[24], sayi2[24], 1'b0, sum[24], carry1[24]);
    full_adder fa_1_26(sayi1[25], sayi2[25], 1'b0, sum[25], carry1[25]);
    full_adder fa_1_27(sayi1[26], sayi2[26], 1'b0, sum[26], carry1[26]);
    full_adder fa_1_28(sayi1[27], sayi2[27], 1'b0, sum[27], carry1[27]);
    full_adder fa_1_29(sayi1[28], sayi2[28], 1'b0, sum[28], carry1[28]);
    full_adder fa_1_30(sayi1[29], sayi2[29], 1'b0, sum[29], carry1[29]);
    full_adder fa_1_31(sayi1[30], sayi2[30], 1'b0, sum[30], carry1[30]);
    full_adder fa_1_32(sayi1[31], sayi2[31], 1'b0, sum[31], carry1[31]);
    full_adder fa_1_33(sayi1[32], sayi2[32], 1'b0, sum[32], carry1[32]);
    full_adder fa_1_34(sayi1[33], sayi2[33], 1'b0, sum[33], carry1[33]);
    full_adder fa_1_35(sayi1[34], sayi2[34], 1'b0, sum[34], carry1[34]);
    full_adder fa_1_36(sayi1[35], sayi2[35], 1'b0, sum[35], carry1[35]);
    full_adder fa_1_37(sayi1[36], sayi2[36], 1'b0, sum[36], carry1[36]);
    full_adder fa_1_38(sayi1[37], sayi2[37], 1'b0, sum[37], carry1[37]);
    full_adder fa_1_39(sayi1[38], sayi2[38], 1'b0, sum[38], carry1[38]);
    full_adder fa_1_40(sayi1[39], sayi2[39], 1'b0, sum[39], carry1[39]);
    full_adder fa_1_41(sayi1[40], sayi2[40], 1'b0, sum[40], carry1[40]);
    full_adder fa_1_42(sayi1[41], sayi2[41], 1'b0, sum[41], carry1[41]);
    full_adder fa_1_43(sayi1[42], sayi2[42], 1'b0, sum[42], carry1[42]);
    full_adder fa_1_44(sayi1[43], sayi2[43], 1'b0, sum[43], carry1[43]);
    full_adder fa_1_45(sayi1[44], sayi2[44], 1'b0, sum[44], carry1[44]);
    full_adder fa_1_46(sayi1[45], sayi2[45], 1'b0, sum[45], carry1[45]);
    full_adder fa_1_47(sayi1[46], sayi2[46], 1'b0, sum[46], carry1[46]);
    full_adder fa_1_48(sayi1[47], sayi2[47], 1'b0, sum[47], carry1[47]);
    full_adder fa_1_49(sayi1[48], sayi2[48], 1'b0, sum[48], carry1[48]);
    full_adder fa_1_50(sayi1[49], sayi2[49], 1'b0, sum[49], carry1[49]);
    full_adder fa_1_51(sayi1[50], sayi2[50], 1'b0, sum[50], carry1[50]);
    full_adder fa_1_52(sayi1[51], sayi2[51], 1'b0, sum[51], carry1[51]);
    full_adder fa_1_53(sayi1[52], sayi2[52], 1'b0, sum[52], carry1[52]);
    full_adder fa_1_54(sayi1[53], sayi2[53], 1'b0, sum[53], carry1[53]);
    full_adder fa_1_55(sayi1[54], sayi2[54], 1'b0, sum[54], carry1[54]);
    full_adder fa_1_56(sayi1[55], sayi2[55], 1'b0, sum[55], carry1[55]);
    full_adder fa_1_57(sayi1[56], sayi2[56], 1'b0, sum[56], carry1[56]);
    full_adder fa_1_58(sayi1[57], sayi2[57], 1'b0, sum[57], carry1[57]);
    full_adder fa_1_59(sayi1[58], sayi2[58], 1'b0, sum[58], carry1[58]);
    full_adder fa_1_60(sayi1[59], sayi2[59], 1'b0, sum[59], carry1[59]);
    full_adder fa_1_61(sayi1[60], sayi2[60], 1'b0, sum[60], carry1[60]);
    full_adder fa_1_62(sayi1[61], sayi2[61], 1'b0, sum[61], carry1[61]);
    full_adder fa_1_63(sayi1[62], sayi2[62], 1'b0, sum[62], carry1[62]);
    full_adder fa_1_64(sayi1[63], sayi2[63], 1'b0, sum[63], carry1[63]);

    full_adder fa_2_1(sum[1], carry1[0], 1'b0, toplam[1], carry2[1]);
    full_adder fa_2_2(sum[2], carry1[1], carry2[1], toplam[2], carry2[2]);
    full_adder fa_2_3(sum[3], carry1[2], carry2[2], toplam[3], carry2[3]);
    full_adder fa_2_4(sum[4], carry1[3], carry2[3], toplam[4], carry2[4]);
    full_adder fa_2_5(sum[5], carry1[4], carry2[4], toplam[5], carry2[5]);
    full_adder fa_2_6(sum[6], carry1[5], carry2[5], toplam[6], carry2[6]);
    full_adder fa_2_7(sum[7], carry1[6], carry2[6], toplam[7], carry2[7]);
    full_adder fa_2_8(sum[8], carry1[7], carry2[7], toplam[8], carry2[8]);
    full_adder fa_2_9(sum[9], carry1[8], carry2[8], toplam[9], carry2[9]);
    full_adder fa_2_10(sum[10], carry1[9], carry2[9], toplam[10], carry2[10]);
    full_adder fa_2_11(sum[11], carry1[10], carry2[10], toplam[11], carry2[11]);
    full_adder fa_2_12(sum[12], carry1[11], carry2[11], toplam[12], carry2[12]);
    full_adder fa_2_13(sum[13], carry1[12], carry2[12], toplam[13], carry2[13]);
    full_adder fa_2_14(sum[14], carry1[13], carry2[13], toplam[14], carry2[14]);
    full_adder fa_2_15(sum[15], carry1[14], carry2[14], toplam[15], carry2[15]);
    full_adder fa_2_16(sum[16], carry1[15], carry2[15], toplam[16], carry2[16]);
    full_adder fa_2_17(sum[17], carry1[16], carry2[16], toplam[17], carry2[17]);
    full_adder fa_2_18(sum[18], carry1[17], carry2[17], toplam[18], carry2[18]);
    full_adder fa_2_19(sum[19], carry1[18], carry2[18], toplam[19], carry2[19]);
    full_adder fa_2_20(sum[20], carry1[19], carry2[19], toplam[20], carry2[20]);
    full_adder fa_2_21(sum[21], carry1[20], carry2[20], toplam[21], carry2[21]);
    full_adder fa_2_22(sum[22], carry1[21], carry2[21], toplam[22], carry2[22]);
    full_adder fa_2_23(sum[23], carry1[22], carry2[22], toplam[23], carry2[23]);
    full_adder fa_2_24(sum[24], carry1[23], carry2[23], toplam[24], carry2[24]);
    full_adder fa_2_25(sum[25], carry1[24], carry2[24], toplam[25], carry2[25]);
    full_adder fa_2_26(sum[26], carry1[25], carry2[25], toplam[26], carry2[26]);
    full_adder fa_2_27(sum[27], carry1[26], carry2[26], toplam[27], carry2[27]);
    full_adder fa_2_28(sum[28], carry1[27], carry2[27], toplam[28], carry2[28]);
    full_adder fa_2_29(sum[29], carry1[28], carry2[28], toplam[29], carry2[29]);
    full_adder fa_2_30(sum[30], carry1[29], carry2[29], toplam[30], carry2[30]);
    full_adder fa_2_31(sum[31], carry1[30], carry2[30], toplam[31], carry2[31]);
    full_adder fa_2_32(sum[32], carry1[31], carry2[31], toplam[32], carry2[32]);
    full_adder fa_2_33(sum[33], carry1[32], carry2[32], toplam[33], carry2[33]);
    full_adder fa_2_34(sum[34], carry1[33], carry2[33], toplam[34], carry2[34]);
    full_adder fa_2_35(sum[35], carry1[34], carry2[34], toplam[35], carry2[35]);
    full_adder fa_2_36(sum[36], carry1[35], carry2[35], toplam[36], carry2[36]);
    full_adder fa_2_37(sum[37], carry1[36], carry2[36], toplam[37], carry2[37]);
    full_adder fa_2_38(sum[38], carry1[37], carry2[37], toplam[38], carry2[38]);
    full_adder fa_2_39(sum[39], carry1[38], carry2[38], toplam[39], carry2[39]);
    full_adder fa_2_40(sum[40], carry1[39], carry2[39], toplam[40], carry2[40]);
    full_adder fa_2_41(sum[41], carry1[40], carry2[40], toplam[41], carry2[41]);
    full_adder fa_2_42(sum[42], carry1[41], carry2[41], toplam[42], carry2[42]);
    full_adder fa_2_43(sum[43], carry1[42], carry2[42], toplam[43], carry2[43]);
    full_adder fa_2_44(sum[44], carry1[43], carry2[43], toplam[44], carry2[44]);
    full_adder fa_2_45(sum[45], carry1[44], carry2[44], toplam[45], carry2[45]);
    full_adder fa_2_46(sum[46], carry1[45], carry2[45], toplam[46], carry2[46]);
    full_adder fa_2_47(sum[47], carry1[46], carry2[46], toplam[47], carry2[47]);
    full_adder fa_2_48(sum[48], carry1[47], carry2[47], toplam[48], carry2[48]);
    full_adder fa_2_49(sum[49], carry1[48], carry2[48], toplam[49], carry2[49]);
    full_adder fa_2_50(sum[50], carry1[49], carry2[49], toplam[50], carry2[50]);
    full_adder fa_2_51(sum[51], carry1[50], carry2[50], toplam[51], carry2[51]);
    full_adder fa_2_52(sum[52], carry1[51], carry2[51], toplam[52], carry2[52]);
    full_adder fa_2_53(sum[53], carry1[52], carry2[52], toplam[53], carry2[53]);
    full_adder fa_2_54(sum[54], carry1[53], carry2[53], toplam[54], carry2[54]);
    full_adder fa_2_55(sum[55], carry1[54], carry2[54], toplam[55], carry2[55]);
    full_adder fa_2_56(sum[56], carry1[55], carry2[55], toplam[56], carry2[56]);
    full_adder fa_2_57(sum[57], carry1[56], carry2[56], toplam[57], carry2[57]);
    full_adder fa_2_58(sum[58], carry1[57], carry2[57], toplam[58], carry2[58]);
    full_adder fa_2_59(sum[59], carry1[58], carry2[58], toplam[59], carry2[59]);
    full_adder fa_2_60(sum[60], carry1[59], carry2[59], toplam[60], carry2[60]);
    full_adder fa_2_61(sum[61], carry1[60], carry2[60], toplam[61], carry2[61]);
    full_adder fa_2_62(sum[62], carry1[61], carry2[61], toplam[62], carry2[62]);
    full_adder fa_2_63(sum[63], carry1[62], carry2[62], toplam[63], carry2[63]);

    assign toplam[0] = sum[0];


endmodule
